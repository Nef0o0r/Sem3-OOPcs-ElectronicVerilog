`timescale 1ns / 1ns

module led_controller_tb();

    reg clk;
    reg [5:0] switches;  // Вход для переключателей
    reg [1:0] buttons;   // Вход для кнопок
    wire [5:0] leds;     // Выход для светодиодов

    // Подключение тестируемого модуля
    led_controller uut (
        .clk(clk),
        .switches(switches),
        .buttons(buttons),
        .leds(leds)
    );

    // Генерация тактового сигнала с периодом 10 нс (частота 100 МГц)
    initial begin
        clk = 0;
        forever #(5) clk = ~clk;
    end

    // Начальные значения для переключателей и кнопок
    initial begin
        switches = 6'b000000; // Все переключатели выключены
        buttons = 6'b000000;  // Все кнопки не нажаты
        
        // Тестовые сценарии
        // Включение всех светодиодов по очереди
        #10 switches[0] = 1;  // Включаем 1-й светодиод
        #10 switches[0] = 0;  // Выключаем

        #10 switches[1] = 1;  // Включаем 2-й светодиод
        #10 switches[1] = 0;  // Выключаем

        #10 switches[2] = 1;  // Включаем 3-й светодиод
        #10 switches[2] = 0;  // Выключаем

        #10 switches[3] = 1;  // Включаем 4-й светодиод
        #10 switches[3] = 0;  // Выключаем

        #10 switches[4] = 1;  // Включаем 5-й светодиод
        #10 switches[4] = 0;  // Выключаем

        #10 switches[5] = 1;  // Включаем 6-й светодиод
        #10 switches[5] = 0;  // Выключаем

        // Инверсия состояния всех светодиодов по очереди
        #10 switches[0] = 1; buttons[0] = 1; // Включаем 1-й и инвертируем
        #10 buttons[0] = 0; // Отпускаем кнопку

        #10 switches[1] = 1; buttons[1] = 1; // Включаем 2-й и инвертируем
        #10 buttons[1] = 0; // Отпускаем кнопку

        #10 switches[2] = 1; buttons[2] = 1; // Включаем 3-й и инвертируем
        #10 buttons[2] = 0; // Отпускаем кнопку

        #10 switches[3] = 1; buttons[3] = 1; // Включаем 4-й и инвертируем
        #10 buttons[3] = 0; // Отпускаем кнопку

        #10 switches[4] = 1; buttons[4] = 1; // Включаем 5-й и инвертируем
        #10 buttons[4] = 0; // Отпускаем кнопку

        #10 switches[5] = 1; buttons[5] = 1; // Включаем 6-й и инвертируем
        #10 buttons[5] = 0; // Отпускаем кнопку
        
        // Завершение симуляции через 200 нс
        #200 $finish;
    end

    // Сохранение результата симуляции в файл VCD
    initial begin
        $dumpfile("led_controller_tb_out.vcd");
        $dumpvars(0, led_controller_tb);
    end

endmodule