`timescale 1ns/1ps

module led_controller_tb;
    reg clk;                  // Тактовый сигнал
    reg [2:0] switches;       // Переключатели
    reg up;                   // Кнопка инверсии
    wire [2:0] leds;          // Светодиоды

    // Экземпляр тестируемого модуля
    led_controller uut (
        .clk(clk),
        .switches(switches),
        .up(up),
        .leds(leds)
    );

    // Генерация тактового сигнала (100 МГц)
    initial begin
        clk = 0;
        forever #5 clk = ~clk; // Период 10 нс
    end

    // Основной блок тестирования
    initial begin
        // Открытие файла для записи результатов
        $dumpfile("led_controller_tb_out.vcd");
        $dumpvars(0, led_controller_tb);

        // Инициализация входов
        switches = 3'b000;
        up = 1;

        // Тест 1: Проверка начального состояния
        #20 switches = 3'b101; // Устанавливаем переключатели
        #20 up = 0;            // Нажимаем кнопку
        #10 up = 1;            // Отпускаем кнопку
        #100;                  // Ждём обработки инверсии

        // Тест 2: Инверсия состояния
        #50 switches = 3'b010; // Изменяем состояние переключателей
        #20 up = 0;            // Нажимаем кнопку для инверсии
        #10 up = 1;            // Отпускаем кнопку
        #100;

        // Тест 3: Включение всех светодиодов
        #50 switches = 3'b111;
        #50;

        // Завершение симуляции
        $finish;
    end
endmodule
