`timescale 1ns / 1ns

module led_controller_tb();

    reg clk;
    reg [2:0] switches;   // Вход для переключателей
    reg [1:0] buttons;    // Вход для кнопок
    wire [5:0] leds;      // Выход для светодиодов

    // Подключение тестируемого модуля
    led_controller uut (
        .clk(clk),
        .switches(switches),
        .buttons(buttons),
        .leds(leds)
    );

    // Генерация тактового сигнала с периодом 10 нс (частота 100 МГц)
    initial begin
        clk = 0;
        forever #(5) clk = ~clk;
    end

    // Начальные значения для переключателей и кнопок
    initial begin
        switches = 3'b000; // Все переключатели выключены
        buttons = 2'b00;   // Кнопки не нажаты

        // Тестовые сценарии
        // Включение светодиодов поочередно с использованием переключателей
        #10 switches[0] = 1;  // Включаем 1-й светодиод
        #10 switches[0] = 0;  // Выключаем 1-й светодиод

        #10 switches[1] = 1;  // Включаем 2-й светодиод
        #10 switches[1] = 0;  // Выключаем 2-й светодиод

        #10 switches[2] = 1;  // Включаем 3-й светодиод
        #10 switches[2] = 0;  // Выключаем 3-й светодиод

        // Включение нескольких светодиодов
        #10 switches = 3'b101;  // Включаем 1-й и 3-й светодиоды
        #10 switches = 3'b010;  // Включаем только 2-й светодиод

        // Инверсия состояния светодиодов
        #10 buttons[0] = 1;  // Нажимаем кнопку для инверсии
        #10 buttons[0] = 0;  // Отпускаем кнопку
        #10 switches = 3'b101; // Проверяем состояние при инверсии

        // Восстановление исходного состояния
        #10 buttons[1] = 1;  // Нажимаем другую кнопку для снятия инверсии
        #10 buttons[1] = 0;  // Отпускаем кнопку

        // Завершение симуляции через 100 нс
        #100 $finish;
    end

    // Сохранение результата симуляции в файл VCD
    initial begin
        $dumpfile("led_controller_tb_out.vcd");
        $dumpvars(0, led_controller_tb);
    end

endmodule